library verilog;
use verilog.vl_types.all;
entity tb_squ_wave is
end tb_squ_wave;
