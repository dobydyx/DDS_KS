module	tb_noise;




endmodule
